module delay_line_2 #(
    parameters
) (
    input clk_inputS
);
    
endmodule